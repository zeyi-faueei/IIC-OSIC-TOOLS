** sch_path: /foss/pdks/sg13g2/libs.tech/xschem/sg13g2_tests/dc_hbt_13g2.sch
**.subckt dc_hbt_13g2
Vce net3 GND 1.5
I0 GND net1 1u
Vc net3 net2 0
.save i(vc)
XQ1 net2 net1 GND GND npn13G2 Nx=1
**** begin user architecture code
.lib cornerHBT.lib hbt_typ
.param temp=27
.control
save all
op
print I(Vc)
reset
dc Vce 0 2 0.01 I0 0 5u 0.1u
write /tmp/test_npn_13G2.raw
quit
.endc
**** end user architecture code
**.ends
.GLOBAL GND
.end
